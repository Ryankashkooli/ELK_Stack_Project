<svg xmlns:xlink="http://www.w3.org/1999/xlink" xmlns="http://www.w3.org/2000/svg" width="1592px" height="530px" viewBox="0 0 1592 530" style="overflow: hidden; display: block; width: 1592px; height: 530px;"><defs/><g style="pointer-events:visiblePainted" transform="translate(2.697163457480727 0)" image-rendering="auto" shape-rendering="auto"><g><path fill="none" stroke="rgb(169,169,169)" d="M 201.66666666666666,240 L 201.66666666666666,250 L 335,250 L 335,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 185,240 L 185,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 168.33333333333334,240 L 168.33333333333334,250 L 35,250 L 35,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 185,140 L 185,180" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 185,60 L 185,80" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 1401.6666666666667,240 L 1401.6666666666667,250 L 1535,250 L 1535,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 1368.3333333333333,240 L 1368.3333333333333,270 L 955,270 L 955,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 1385,240 L 1385,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 955,140 L 955,150 L 1385,150 L 1385,180" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 1072.5,240 L 1072.5,260 L 945,260 L 945,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 1097.5,240 L 1097.5,250 L 1235,250 L 1235,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 945,140 L 945,160 L 1085,160 L 1085,180" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 951.6666666666666,240 L 951.6666666666666,250 L 1085,250 L 1085,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 647.5,440 L 647.5,470" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 622.5,440 L 622.5,450 L 497.5,450 L 497.5,470" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 635,360 L 635,380" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 918.3333333333334,240 L 918.3333333333334,260 L 651.6666666666666,260 L 651.6666666666666,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 935,240 L 935,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 935,140 L 935,180" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 785,240 L 785,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 768.3333333333334,240 L 768.3333333333334,250 L 635,250 L 635,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 801.6666666666666,240 L 801.6666666666666,270 L 925,270 L 925,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 925,140 L 925,160 L 785,160 L 785,180" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 601.6666666666667,240 L 601.6666666666667,250 L 485,250 L 485,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 618.3333333333334,240 L 618.3333333333334,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 635,240 L 635,280 L 915,280 L 915,300" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 915,140 L 915,150 L 618.3333333333334,150 L 618.3333333333334,180" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 935,60 L 935,80" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 210,30 L 910,30" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g><path fill="none" stroke="rgb(169,169,169)" d="M 910,30 L 210,30" stroke-opacity="1" stroke-width="1" stroke-linecap="butt" stroke-linejoin="miter" stroke-miterlimit="10"/></g><g transform="translate(160 0)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_0" x1="9.88" y1="8.59" x2="11.52" y2="10.23" gradientTransform="rotate(-.08 -285.464 -1454.08)" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#86d633"/><stop offset=".24" stop-color="#83d232"/><stop offset=".5" stop-color="#7cc52f"/><stop offset=".76" stop-color="#6fb02a"/><stop offset="1" stop-color="#5e9624"/></linearGradient><linearGradient id="ygc3_1" x1="6.18" y1="8.59" x2="7.81" y2="10.23"/><linearGradient id="ygc3_2" x1="2.48" y1="8.59" x2="4.11" y2="10.23"/></defs><title>Icon-networking-61</title><circle cx="12.74" cy="8.99" r="1.16" fill="url(#ygc3_0)"/><circle cx="9.04" cy="9" r="1.16" fill="url(#ygc3_1)"/><circle cx="5.34" cy="9" r="1.16" fill="url(#ygc3_2)"/><path d="M6.182 13.638l-.664.665a.3.3 0 0 1-.424 0L.18 9.404a.6.6 0 0 1-.001-.848l.663-.666 5.34 5.324a.3.3 0 0 1 0 .425z" fill="#50e6ff"/><path d="M5.418 3.708l.666.664a.3.3 0 0 1 0 .424L.838 10.057l-.666-.663a.6.6 0 0 1-.001-.849L4.994 3.71a.3.3 0 0 1 .424 0z" fill="#1490df"/><path d="M17.157 7.88l.663.666a.6.6 0 0 1 0 .848l-4.915 4.9a.3.3 0 0 1-.424 0l-.664-.666a.3.3 0 0 1 0-.424l5.34-5.324z" fill="#50e6ff"/><path d="M17.818 9.387l-.665.664-5.247-5.261a.3.3 0 0 1 0-.425l.674-.67a.3.3 0 0 1 .424 0l4.823 4.836a.6.6 0 0 1-.002.849z" fill="#1490df"/></g></svg>
        </g></g><g transform="translate(160 80)"><g transform="scale(1.0)">
            <svg svgBox="0 0 50 50" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><path d="M49.7 25.7c.5-.5.4-1.3 0-1.8l-2.4-2.4L36.5 11c-.5-.5-1.2-.5-1.7 0s-.6 1.3 0 1.8l11.3 11.1c.5.5.5 1.3 0 1.8L34.6 37.2c-.5.5-.5 1.3 0 1.8s1.3.4 1.7 0L47 28.4l.1-.1 2.6-2.6zm-49.4 0c-.5-.5-.4-1.3 0-1.8l2.4-2.4L13.5 11c.5-.5 1.2-.5 1.7 0s.6 1.3 0 1.8L4.1 23.9c-.5.5-.5 1.3 0 1.8l11.3 11.5c.5.5.5 1.3 0 1.8s-1.3.4-1.7 0L2.8 28.5l-.1-.1-2.4-2.7z" fill="#3999C6"/><path d="M28.4 24.8c0 1.9-1.6 3.3-3.3 3.3-1.7 0-3.5-1.6-3.5-3.3s1.4-3.3 3.5-3.3c2 0 3.3 1.6 3.3 3.3z" fill="#7fba00"/></g></svg>
        </g></g><g transform="translate(160 180)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_3" x1="9.01" y1="16.5" x2="9.01" y2="1.5" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#5e9641"/><stop offset=".34" stop-color="#6baa42"/><stop offset=".67" stop-color="#73b743"/><stop offset="1" stop-color="#76bb43"/></linearGradient></defs><title>Icon-networking-80</title><path d="M15.89 2.91h1.27a.34.34 0 0 1 .34.34v3.5a.34.34 0 0 1-.34.34h-1.27V2.91zm0 6.09h1.27a.34.34 0 0 1 .34.34v5.86a.34.34 0 0 1-.34.34h-1.27V9z" fill="#ffca00"/><rect x="2.13" y="1.5" width="13.76" height="15" rx=".69" fill="url(#ygc3_3)"/><path d="M5.9 12.9h-.71a.2.2 0 0 1-.19-.21V4.34a.19.19 0 0 1 .19-.2h1.93a.19.19 0 0 1 .19.2.2.2 0 0 1-.19.21H5.38v7.93h.52a.2.2 0 0 1 .19.21.21.21 0 0 1-.19.21z" fill="#b4ec36"/><path d="M6 13.92H4.4a.2.2 0 0 1-.19-.21L4.08 3.38a.2.2 0 0 1 .06-.15.16.16 0 0 1 .13-.06h2.85v.41H4.47l.12 9.92H6zm6-.92h-1.59a.19.19 0 0 1-.14-.07.18.18 0 0 1-.06-.14V7.9a.19.19 0 0 1 .19-.2h.91V5.45h.38v2.44a.2.2 0 0 1-.18.21h-.91v4.42H12z" fill="#b4ec36"/><rect x="7.07" y="2.29" width="6.14" height="3.11" rx=".26" fill="#365615"/><rect x="5.86" y="12.69" width="4.9" height="1.09" rx=".26" transform="rotate(90 8.305 13.235)" fill="#365615"/><rect x="3.99" y="12.71" width="4.9" height="1.09" rx=".26" transform="rotate(90 6.44 13.26)" fill="#365615"/><rect x="9.98" y="12.71" width="4.9" height="1.09" rx=".26" transform="rotate(90 12.425 13.255)" fill="#f2f2f2"/><ellipse cx="8.11" cy="8.06" rx="1.04" ry="1.12" fill="#f2f2f2"/><path d="M2.11 12.25H.84a.34.34 0 0 1-.34-.3V6.09a.34.34 0 0 1 .34-.34h1.27v6.5z" fill="#3b3b3b"/></g></svg>
        </g></g><g transform="translate(310 300)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_4" x1="8.88" y1="12.21" x2="8.88" y2=".21" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#0078d4"/><stop offset=".82" stop-color="#5ea0ef"/></linearGradient><linearGradient id="ygc3_5" x1="8.88" y1="16.84" x2="8.88" y2="12.21" gradientUnits="userSpaceOnUse"><stop offset=".15" stop-color="#ccc"/><stop offset="1" stop-color="#707070"/></linearGradient></defs><title>Icon-compute-21</title><rect x="-.12" y=".21" width="18" height="12" rx=".6" fill="url(#ygc3_4)"/><path fill="#50e6ff" d="M11.88 4.46v3.49l-3 1.76v-3.5l3-1.75z"/><path fill="#c3f1ff" d="M11.88 4.46l-3 1.76-3-1.76 3-1.75 3 1.75z"/><path fill="#9cebff" d="M8.88 6.22v3.49l-3-1.76V4.46l3 1.76z"/><path fill="#c3f1ff" d="M5.88 7.95l3-1.74v3.5l-3-1.76z"/><path fill="#9cebff" d="M11.88 7.95l-3-1.74v3.5l3-1.76z"/><path d="M12.49 15.84c-1.78-.28-1.85-1.56-1.85-3.63H7.11c0 2.07-.06 3.35-1.84 3.63a1 1 0 0 0-.89 1h9a1 1 0 0 0-.89-1z" fill="url(#ygc3_5)"/></g></svg>
        </g></g><g transform="translate(160 300)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_6" x1="9.01" y1=".75" x2="9.01" y2="17.25" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#5ea0ef"/><stop offset=".18" stop-color="#559cec"/><stop offset=".47" stop-color="#3c91e5"/><stop offset=".84" stop-color="#1380da"/><stop offset="1" stop-color="#0078d4"/></linearGradient></defs><title>Icon-networking-67</title><path d="M16.36 8.4c0 4.84-5.85 8.74-7.12 9.53a.46.46 0 0 1-.48 0c-1.27-.79-7.12-4.69-7.12-9.53V2.58a.46.46 0 0 1 .45-.46C6.64 2 5.59 0 9 0s2.36 2 6.91 2.12a.46.46 0 0 1 .45.46z" fill="#0078d4"/><path d="M15.75 8.45c0 4.44-5.36 8-6.53 8.74a.43.43 0 0 1-.44 0c-1.17-.72-6.53-4.3-6.53-8.74V3.11a.42.42 0 0 1 .41-.42C6.83 2.58 5.87.75 9 .75s2.17 1.83 6.34 1.94a.42.42 0 0 1 .41.42z" fill="#6bb9f2"/><path d="M9 9V.75c3.13 0 2.17 1.83 6.34 1.94a.43.43 0 0 1 .41.43v5.34a4.89 4.89 0 0 1 0 .54zm0 0H2.28c.4 4.18 5.38 7.5 6.5 8.19a.39.39 0 0 0 .18.06H9z" fill="url(#ygc3_6)"/><path d="M2.66 2.69C6.83 2.58 5.87.75 9 .75V9H2.28a4.89 4.89 0 0 1 0-.54V3.12a.43.43 0 0 1 .38-.43zM15.72 9H9v8.25a.39.39 0 0 0 .18-.06c1.16-.69 6.14-4.01 6.54-8.19z" fill="#50e6ff"/></g></svg>
        </g></g><g transform="translate(10 300)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_7" x1="9" y1="15.83" x2="9" y2="5.79" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#32bedd"/><stop offset=".18" stop-color="#32caea"/><stop offset=".41" stop-color="#32d2f2"/><stop offset=".78" stop-color="#32d4f5"/></linearGradient></defs><title>Icon-networking-69</title><path d="M.5 5.79h17v9.48a.57.57 0 0 1-.57.57H1.07a.57.57 0 0 1-.57-.57V5.79z" fill="url(#ygc3_7)"/><path d="M1.07 2.17h15.86a.57.57 0 0 1 .57.57v3.05H.5V2.73a.57.57 0 0 1 .57-.56z" fill="#767676"/><circle cx="12.82" cy="10.19" r="1.38" fill="#f2f2f2"/><circle cx="9.06" cy="10.19" r="1.38" fill="#f2f2f2"/><circle cx="5.18" cy="10.19" r="1.38" fill="#f2f2f2"/><rect x="2.79" y="3.25" width="12.43" height="1.46" rx=".28" fill="#f2f2f2"/></g></svg>
        </g></g><g transform="translate(910 0)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_8" x1="9.88" y1="8.59" x2="11.52" y2="10.23" gradientTransform="rotate(-.08 -285.464 -1454.08)" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#86d633"/><stop offset=".24" stop-color="#83d232"/><stop offset=".5" stop-color="#7cc52f"/><stop offset=".76" stop-color="#6fb02a"/><stop offset="1" stop-color="#5e9624"/></linearGradient><linearGradient id="ygc3_9" x1="6.18" y1="8.59" x2="7.81" y2="10.23"/><linearGradient id="ygc3_10" x1="2.48" y1="8.59" x2="4.11" y2="10.23"/></defs><title>Icon-networking-61</title><circle cx="12.74" cy="8.99" r="1.16" fill="url(#ygc3_8)"/><circle cx="9.04" cy="9" r="1.16" fill="url(#ygc3_9)"/><circle cx="5.34" cy="9" r="1.16" fill="url(#ygc3_10)"/><path d="M6.182 13.638l-.664.665a.3.3 0 0 1-.424 0L.18 9.404a.6.6 0 0 1-.001-.848l.663-.666 5.34 5.324a.3.3 0 0 1 0 .425z" fill="#50e6ff"/><path d="M5.418 3.708l.666.664a.3.3 0 0 1 0 .424L.838 10.057l-.666-.663a.6.6 0 0 1-.001-.849L4.994 3.71a.3.3 0 0 1 .424 0z" fill="#1490df"/><path d="M17.157 7.88l.663.666a.6.6 0 0 1 0 .848l-4.915 4.9a.3.3 0 0 1-.424 0l-.664-.666a.3.3 0 0 1 0-.424l5.34-5.324z" fill="#50e6ff"/><path d="M17.818 9.387l-.665.664-5.247-5.261a.3.3 0 0 1 0-.425l.674-.67a.3.3 0 0 1 .424 0l4.823 4.836a.6.6 0 0 1-.002.849z" fill="#1490df"/></g></svg>
        </g></g><g transform="translate(910 80)"><g transform="scale(1.0)">
            <svg svgBox="0 0 50 50" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><path d="M49.7 25.7c.5-.5.4-1.3 0-1.8l-2.4-2.4L36.5 11c-.5-.5-1.2-.5-1.7 0s-.6 1.3 0 1.8l11.3 11.1c.5.5.5 1.3 0 1.8L34.6 37.2c-.5.5-.5 1.3 0 1.8s1.3.4 1.7 0L47 28.4l.1-.1 2.6-2.6zm-49.4 0c-.5-.5-.4-1.3 0-1.8l2.4-2.4L13.5 11c.5-.5 1.2-.5 1.7 0s.6 1.3 0 1.8L4.1 23.9c-.5.5-.5 1.3 0 1.8l11.3 11.5c.5.5.5 1.3 0 1.8s-1.3.4-1.7 0L2.8 28.5l-.1-.1-2.4-2.7z" fill="#3999C6"/><path d="M28.4 24.8c0 1.9-1.6 3.3-3.3 3.3-1.7 0-3.5-1.6-3.5-3.3s1.4-3.3 3.5-3.3c2 0 3.3 1.6 3.3 3.3z" fill="#7fba00"/></g></svg>
        </g></g><g transform="translate(1360 180)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_11" x1="9.01" y1="16.5" x2="9.01" y2="1.5" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#5e9641"/><stop offset=".34" stop-color="#6baa42"/><stop offset=".67" stop-color="#73b743"/><stop offset="1" stop-color="#76bb43"/></linearGradient></defs><title>Icon-networking-80</title><path d="M15.89 2.91h1.27a.34.34 0 0 1 .34.34v3.5a.34.34 0 0 1-.34.34h-1.27V2.91zm0 6.09h1.27a.34.34 0 0 1 .34.34v5.86a.34.34 0 0 1-.34.34h-1.27V9z" fill="#ffca00"/><rect x="2.13" y="1.5" width="13.76" height="15" rx=".69" fill="url(#ygc3_11)"/><path d="M5.9 12.9h-.71a.2.2 0 0 1-.19-.21V4.34a.19.19 0 0 1 .19-.2h1.93a.19.19 0 0 1 .19.2.2.2 0 0 1-.19.21H5.38v7.93h.52a.2.2 0 0 1 .19.21.21.21 0 0 1-.19.21z" fill="#b4ec36"/><path d="M6 13.92H4.4a.2.2 0 0 1-.19-.21L4.08 3.38a.2.2 0 0 1 .06-.15.16.16 0 0 1 .13-.06h2.85v.41H4.47l.12 9.92H6zm6-.92h-1.59a.19.19 0 0 1-.14-.07.18.18 0 0 1-.06-.14V7.9a.19.19 0 0 1 .19-.2h.91V5.45h.38v2.44a.2.2 0 0 1-.18.21h-.91v4.42H12z" fill="#b4ec36"/><rect x="7.07" y="2.29" width="6.14" height="3.11" rx=".26" fill="#365615"/><rect x="5.86" y="12.69" width="4.9" height="1.09" rx=".26" transform="rotate(90 8.305 13.235)" fill="#365615"/><rect x="3.99" y="12.71" width="4.9" height="1.09" rx=".26" transform="rotate(90 6.44 13.26)" fill="#365615"/><rect x="9.98" y="12.71" width="4.9" height="1.09" rx=".26" transform="rotate(90 12.425 13.255)" fill="#f2f2f2"/><ellipse cx="8.11" cy="8.06" rx="1.04" ry="1.12" fill="#f2f2f2"/><path d="M2.11 12.25H.84a.34.34 0 0 1-.34-.3V6.09a.34.34 0 0 1 .34-.34h1.27v6.5z" fill="#3b3b3b"/></g></svg>
        </g></g><g transform="translate(1510 300)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_12" x1="8.88" y1="12.21" x2="8.88" y2=".21" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#0078d4"/><stop offset=".82" stop-color="#5ea0ef"/></linearGradient><linearGradient id="ygc3_13" x1="8.88" y1="16.84" x2="8.88" y2="12.21" gradientUnits="userSpaceOnUse"><stop offset=".15" stop-color="#ccc"/><stop offset="1" stop-color="#707070"/></linearGradient></defs><title>Icon-compute-21</title><rect x="-.12" y=".21" width="18" height="12" rx=".6" fill="url(#ygc3_12)"/><path fill="#50e6ff" d="M11.88 4.46v3.49l-3 1.76v-3.5l3-1.75z"/><path fill="#c3f1ff" d="M11.88 4.46l-3 1.76-3-1.76 3-1.75 3 1.75z"/><path fill="#9cebff" d="M8.88 6.22v3.49l-3-1.76V4.46l3 1.76z"/><path fill="#c3f1ff" d="M5.88 7.95l3-1.74v3.5l-3-1.76z"/><path fill="#9cebff" d="M11.88 7.95l-3-1.74v3.5l3-1.76z"/><path d="M12.49 15.84c-1.78-.28-1.85-1.56-1.85-3.63H7.11c0 2.07-.06 3.35-1.84 3.63a1 1 0 0 0-.89 1h9a1 1 0 0 0-.89-1z" fill="url(#ygc3_13)"/></g></svg>
        </g></g><g transform="translate(910 300)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_14" x1="9.01" y1=".75" x2="9.01" y2="17.25" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#5ea0ef"/><stop offset=".18" stop-color="#559cec"/><stop offset=".47" stop-color="#3c91e5"/><stop offset=".84" stop-color="#1380da"/><stop offset="1" stop-color="#0078d4"/></linearGradient></defs><title>Icon-networking-67</title><path d="M16.36 8.4c0 4.84-5.85 8.74-7.12 9.53a.46.46 0 0 1-.48 0c-1.27-.79-7.12-4.69-7.12-9.53V2.58a.46.46 0 0 1 .45-.46C6.64 2 5.59 0 9 0s2.36 2 6.91 2.12a.46.46 0 0 1 .45.46z" fill="#0078d4"/><path d="M15.75 8.45c0 4.44-5.36 8-6.53 8.74a.43.43 0 0 1-.44 0c-1.17-.72-6.53-4.3-6.53-8.74V3.11a.42.42 0 0 1 .41-.42C6.83 2.58 5.87.75 9 .75s2.17 1.83 6.34 1.94a.42.42 0 0 1 .41.42z" fill="#6bb9f2"/><path d="M9 9V.75c3.13 0 2.17 1.83 6.34 1.94a.43.43 0 0 1 .41.43v5.34a4.89 4.89 0 0 1 0 .54zm0 0H2.28c.4 4.18 5.38 7.5 6.5 8.19a.39.39 0 0 0 .18.06H9z" fill="url(#ygc3_14)"/><path d="M2.66 2.69C6.83 2.58 5.87.75 9 .75V9H2.28a4.89 4.89 0 0 1 0-.54V3.12a.43.43 0 0 1 .38-.43zM15.72 9H9v8.25a.39.39 0 0 0 .18-.06c1.16-.69 6.14-4.01 6.54-8.19z" fill="#50e6ff"/></g></svg>
        </g></g><g transform="translate(1360 300)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_15" x1="9" y1="15.83" x2="9" y2="5.79" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#32bedd"/><stop offset=".18" stop-color="#32caea"/><stop offset=".41" stop-color="#32d2f2"/><stop offset=".78" stop-color="#32d4f5"/></linearGradient></defs><title>Icon-networking-69</title><path d="M.5 5.79h17v9.48a.57.57 0 0 1-.57.57H1.07a.57.57 0 0 1-.57-.57V5.79z" fill="url(#ygc3_15)"/><path d="M1.07 2.17h15.86a.57.57 0 0 1 .57.57v3.05H.5V2.73a.57.57 0 0 1 .57-.56z" fill="#767676"/><circle cx="12.82" cy="10.19" r="1.38" fill="#f2f2f2"/><circle cx="9.06" cy="10.19" r="1.38" fill="#f2f2f2"/><circle cx="5.18" cy="10.19" r="1.38" fill="#f2f2f2"/><rect x="2.79" y="3.25" width="12.43" height="1.46" rx=".28" fill="#f2f2f2"/></g></svg>
        </g></g><g transform="translate(1060 180)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_16" x1="9.01" y1="16.5" x2="9.01" y2="1.5" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#5e9641"/><stop offset=".34" stop-color="#6baa42"/><stop offset=".67" stop-color="#73b743"/><stop offset="1" stop-color="#76bb43"/></linearGradient></defs><title>Icon-networking-80</title><path d="M15.89 2.91h1.27a.34.34 0 0 1 .34.34v3.5a.34.34 0 0 1-.34.34h-1.27V2.91zm0 6.09h1.27a.34.34 0 0 1 .34.34v5.86a.34.34 0 0 1-.34.34h-1.27V9z" fill="#ffca00"/><rect x="2.13" y="1.5" width="13.76" height="15" rx=".69" fill="url(#ygc3_16)"/><path d="M5.9 12.9h-.71a.2.2 0 0 1-.19-.21V4.34a.19.19 0 0 1 .19-.2h1.93a.19.19 0 0 1 .19.2.2.2 0 0 1-.19.21H5.38v7.93h.52a.2.2 0 0 1 .19.21.21.21 0 0 1-.19.21z" fill="#b4ec36"/><path d="M6 13.92H4.4a.2.2 0 0 1-.19-.21L4.08 3.38a.2.2 0 0 1 .06-.15.16.16 0 0 1 .13-.06h2.85v.41H4.47l.12 9.92H6zm6-.92h-1.59a.19.19 0 0 1-.14-.07.18.18 0 0 1-.06-.14V7.9a.19.19 0 0 1 .19-.2h.91V5.45h.38v2.44a.2.2 0 0 1-.18.21h-.91v4.42H12z" fill="#b4ec36"/><rect x="7.07" y="2.29" width="6.14" height="3.11" rx=".26" fill="#365615"/><rect x="5.86" y="12.69" width="4.9" height="1.09" rx=".26" transform="rotate(90 8.305 13.235)" fill="#365615"/><rect x="3.99" y="12.71" width="4.9" height="1.09" rx=".26" transform="rotate(90 6.44 13.26)" fill="#365615"/><rect x="9.98" y="12.71" width="4.9" height="1.09" rx=".26" transform="rotate(90 12.425 13.255)" fill="#f2f2f2"/><ellipse cx="8.11" cy="8.06" rx="1.04" ry="1.12" fill="#f2f2f2"/><path d="M2.11 12.25H.84a.34.34 0 0 1-.34-.3V6.09a.34.34 0 0 1 .34-.34h1.27v6.5z" fill="#3b3b3b"/></g></svg>
        </g></g><g transform="translate(1210 300)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_17" x1="9" y1="15.83" x2="9" y2="5.79" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#32bedd"/><stop offset=".18" stop-color="#32caea"/><stop offset=".41" stop-color="#32d2f2"/><stop offset=".78" stop-color="#32d4f5"/></linearGradient></defs><title>Icon-networking-69</title><path d="M.5 5.79h17v9.48a.57.57 0 0 1-.57.57H1.07a.57.57 0 0 1-.57-.57V5.79z" fill="url(#ygc3_17)"/><path d="M1.07 2.17h15.86a.57.57 0 0 1 .57.57v3.05H.5V2.73a.57.57 0 0 1 .57-.56z" fill="#767676"/><circle cx="12.82" cy="10.19" r="1.38" fill="#f2f2f2"/><circle cx="9.06" cy="10.19" r="1.38" fill="#f2f2f2"/><circle cx="5.18" cy="10.19" r="1.38" fill="#f2f2f2"/><rect x="2.79" y="3.25" width="12.43" height="1.46" rx=".28" fill="#f2f2f2"/></g></svg>
        </g></g><g transform="translate(910 180)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_18" x1="9.01" y1="16.5" x2="9.01" y2="1.5" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#5e9641"/><stop offset=".34" stop-color="#6baa42"/><stop offset=".67" stop-color="#73b743"/><stop offset="1" stop-color="#76bb43"/></linearGradient></defs><title>Icon-networking-80</title><path d="M15.89 2.91h1.27a.34.34 0 0 1 .34.34v3.5a.34.34 0 0 1-.34.34h-1.27V2.91zm0 6.09h1.27a.34.34 0 0 1 .34.34v5.86a.34.34 0 0 1-.34.34h-1.27V9z" fill="#ffca00"/><rect x="2.13" y="1.5" width="13.76" height="15" rx=".69" fill="url(#ygc3_18)"/><path d="M5.9 12.9h-.71a.2.2 0 0 1-.19-.21V4.34a.19.19 0 0 1 .19-.2h1.93a.19.19 0 0 1 .19.2.2.2 0 0 1-.19.21H5.38v7.93h.52a.2.2 0 0 1 .19.21.21.21 0 0 1-.19.21z" fill="#b4ec36"/><path d="M6 13.92H4.4a.2.2 0 0 1-.19-.21L4.08 3.38a.2.2 0 0 1 .06-.15.16.16 0 0 1 .13-.06h2.85v.41H4.47l.12 9.92H6zm6-.92h-1.59a.19.19 0 0 1-.14-.07.18.18 0 0 1-.06-.14V7.9a.19.19 0 0 1 .19-.2h.91V5.45h.38v2.44a.2.2 0 0 1-.18.21h-.91v4.42H12z" fill="#b4ec36"/><rect x="7.07" y="2.29" width="6.14" height="3.11" rx=".26" fill="#365615"/><rect x="5.86" y="12.69" width="4.9" height="1.09" rx=".26" transform="rotate(90 8.305 13.235)" fill="#365615"/><rect x="3.99" y="12.71" width="4.9" height="1.09" rx=".26" transform="rotate(90 6.44 13.26)" fill="#365615"/><rect x="9.98" y="12.71" width="4.9" height="1.09" rx=".26" transform="rotate(90 12.425 13.255)" fill="#f2f2f2"/><ellipse cx="8.11" cy="8.06" rx="1.04" ry="1.12" fill="#f2f2f2"/><path d="M2.11 12.25H.84a.34.34 0 0 1-.34-.3V6.09a.34.34 0 0 1 .34-.34h1.27v6.5z" fill="#3b3b3b"/></g></svg>
        </g></g><g transform="translate(1060 300)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_19" x1="8.88" y1="12.21" x2="8.88" y2=".21" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#0078d4"/><stop offset=".82" stop-color="#5ea0ef"/></linearGradient><linearGradient id="ygc3_20" x1="8.88" y1="16.84" x2="8.88" y2="12.21" gradientUnits="userSpaceOnUse"><stop offset=".15" stop-color="#ccc"/><stop offset="1" stop-color="#707070"/></linearGradient></defs><title>Icon-compute-21</title><rect x="-.12" y=".21" width="18" height="12" rx=".6" fill="url(#ygc3_19)"/><path fill="#50e6ff" d="M11.88 4.46v3.49l-3 1.76v-3.5l3-1.75z"/><path fill="#c3f1ff" d="M11.88 4.46l-3 1.76-3-1.76 3-1.75 3 1.75z"/><path fill="#9cebff" d="M8.88 6.22v3.49l-3-1.76V4.46l3 1.76z"/><path fill="#c3f1ff" d="M5.88 7.95l3-1.74v3.5l-3-1.76z"/><path fill="#9cebff" d="M11.88 7.95l-3-1.74v3.5l3-1.76z"/><path d="M12.49 15.84c-1.78-.28-1.85-1.56-1.85-3.63H7.11c0 2.07-.06 3.35-1.84 3.63a1 1 0 0 0-.89 1h9a1 1 0 0 0-.89-1z" fill="url(#ygc3_20)"/></g></svg>
        </g></g><g transform="translate(610 300)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_21" x1="10.31" y1="12.7" x2="10.31" y2="6.83" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#0078d4"/><stop offset=".82" stop-color="#5ea0ef"/></linearGradient><linearGradient id="ygc3_22" x1="10.31" y1="14.97" x2="10.31" y2="12.7" gradientUnits="userSpaceOnUse"><stop offset=".15" stop-color="#ccc"/><stop offset="1" stop-color="#707070"/></linearGradient></defs><title>Icon-compute-25</title><path fill="#0078d4" d="M2.12.5h1.97v.57H2.12zm14.51.57h.32v.31h.55V.5h-.87v.57zM1.41 16.89h-.28v-.32H.5v.93h.91v-.61zm15.54-.29v.29h-.32v.61h.87v-.9h-.55zM1.13 1.36v-.29h.28V.5H.5v.86h.63z"/><rect x="3.37" y="3.55" width="8.79" height="5.88" rx=".29" fill="#0078d4"/><path fill="#50e6ff" d="M9.23 5.64v1.71l-1.46.86V6.49l1.46-.85z"/><path fill="#c3f1ff" d="M9.23 5.64l-1.46.86-1.47-.86 1.47-.86 1.46.86z"/><path fill="#9cebff" d="M7.77 6.5v1.71L6.3 7.35V5.64l1.47.86z"/><rect x="5.91" y="6.83" width="8.79" height="5.88" rx=".29" fill="url(#ygc3_21)"/><path fill="#50e6ff" d="M11.77 8.91v1.71l-1.46.86V9.77l1.46-.86z"/><path fill="#c3f1ff" d="M11.77 8.91l-1.46.86-1.47-.86 1.47-.86 1.46.86z"/><path fill="#9cebff" d="M10.31 9.77v1.71l-1.47-.86V8.91l1.47.86z"/><path fill="#c3f1ff" d="M8.84 10.62l1.47-.85v1.71l-1.47-.86z"/><path fill="#9cebff" d="M11.77 10.62l-1.46-.85v1.71l1.46-.86z"/><path d="M12.07 14.48c-.87-.14-.9-.77-.9-1.78H9.44c0 1 0 1.64-.9 1.78a.51.51 0 0 0-.43.49h4.4a.51.51 0 0 0-.44-.49z" fill="url(#ygc3_22)"/><path fill="#0078d4" d="M5.07.5h1.97v.57H5.07zm2.94 0h1.97v.57H8.01zm2.95 0h1.97v.57h-1.97zm2.95 0h1.97v.57h-1.97zM2.14 16.89h1.97v.57H2.14zm2.94 0h1.97v.57H5.08zm2.95 0H10v.57H8.03zm2.95 0h1.97v.57h-1.97zm2.94 0h1.97v.57h-1.97zm3.01-14.84h.57v1.97h-.57zm0 2.94h.57v1.97h-.57zm0 2.95h.57v1.97h-.57zm0 2.94h.57v1.97h-.57zm0 2.95h.57v1.97h-.57zM.5 2.03h.57V4H.5zm0 2.95h.57v1.97H.5zm0 2.94h.57v1.97H.5zm0 2.95h.57v1.97H.5zm0 2.94h.57v1.97H.5z"/></g></svg>
        </g></g><g transform="translate(610 380)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_23" x1="9" y1="19.85" x2="9" y2="-1.02" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#5e9624"/><stop offset=".02" stop-color="#5f9724"/><stop offset="1" stop-color="#76bc2d"/></linearGradient></defs><title>Icon-networking-62</title><path d="M.18 8.57L8.57.18a.6.6 0 0 1 .86 0l8.39 8.39a.6.6 0 0 1 0 .86l-8.4 8.4a.6.6 0 0 1-.84 0l-8.4-8.4a.6.6 0 0 1 0-.86z" fill="url(#ygc3_23)"/><path d="M11.2 4L9.08 1.89a.12.12 0 0 0-.16 0L6.8 4a.1.1 0 0 0 .08.18h1.24a.11.11 0 0 1 .11.11v2a.11.11 0 0 0 .11.11h1.32a.11.11 0 0 0 .11-.11v-2a.11.11 0 0 1 .11-.11h1.24A.1.1 0 0 0 11.2 4zM4 6.61L1.9 8.74a.11.11 0 0 0 0 .15L4 11a.11.11 0 0 0 .19-.08V9.69a.11.11 0 0 1 .11-.11h2a.1.1 0 0 0 .1-.11V8.15A.1.1 0 0 0 6.33 8h-2a.1.1 0 0 1-.11-.1V6.69A.11.11 0 0 0 4 6.61zM14.08 11l2.13-2.12a.11.11 0 0 0 0-.15l-2.13-2.12a.11.11 0 0 0-.18.08v1.25a.1.1 0 0 1-.11.1h-2a.1.1 0 0 0-.1.11v1.32a.1.1 0 0 0 .1.11h2a.11.11 0 0 1 .11.11v1.24a.11.11 0 0 0 .18.07z" fill="#b4ec36"/><path d="M11.79 9a2.79 2.79 0 1 0-3.54 2.67v.95a1.71 1.71 0 1 0 1.57 0v-1A2.77 2.77 0 0 0 11.79 9z" fill="#fff"/><circle cx="9.01" cy="8.99" r="1.62" fill="#5ea0ef"/></g></svg>
        </g></g><g transform="translate(622.5 470)"><g transform="scale(1.0)">
            <svg svgBox="0 0 50 50" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><polygon points="27.1,21.8 22.9,21.8 19.7,50 30.3,50" fill="#59b4d9"/><path d="M40.3 22.5C40.3 14 33.5 7.1 25 7.1S9.7 14 9.7 22.5c0 5.6 3 10.5 7.6 13.2.5-.8.9-1.6 1.3-2.3-3.7-2.2-6.2-6.2-6.2-10.9 0-7 5.7-12.7 12.7-12.7 7 0 12.7 5.7 12.7 12.7 0 4.6-2.5 8.7-6.2 10.9.4.7.9 1.5 1.3 2.3 4.4-2.7 7.4-7.6 7.4-13.2" opacity=".5" fill="#3e3e3e"/><path d="M13.7 41.9c.4-.8.9-1.6 1.3-2.4-5.9-3.4-9.8-9.8-9.8-17.1C5.2 11.6 14.1 2.7 25 2.7s19.8 8.9 19.8 19.8c0 7.3-4 13.6-9.8 17.1.4.8.9 1.6 1.3 2.4 6.7-3.9 11.2-11.1 11.2-19.4C47.5 10.1 37.4 0 25 0S2.5 10.1 2.5 22.5c0 8.2 4.6 15.5 11.2 19.4" opacity=".2" fill="#3e3e3e"/><circle cx="25" cy="22.6" r="6.8" fill="#0072c6"/></g></svg>
        </g></g><g transform="translate(472.5 470)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_24" x1="9" y1="15.83" x2="9" y2="5.79" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#32bedd"/><stop offset=".18" stop-color="#32caea"/><stop offset=".41" stop-color="#32d2f2"/><stop offset=".78" stop-color="#32d4f5"/></linearGradient></defs><title>Icon-networking-69</title><path d="M.5 5.79h17v9.48a.57.57 0 0 1-.57.57H1.07a.57.57 0 0 1-.57-.57V5.79z" fill="url(#ygc3_24)"/><path d="M1.07 2.17h15.86a.57.57 0 0 1 .57.57v3.05H.5V2.73a.57.57 0 0 1 .57-.56z" fill="#767676"/><circle cx="12.82" cy="10.19" r="1.38" fill="#f2f2f2"/><circle cx="9.06" cy="10.19" r="1.38" fill="#f2f2f2"/><circle cx="5.18" cy="10.19" r="1.38" fill="#f2f2f2"/><rect x="2.79" y="3.25" width="12.43" height="1.46" rx=".28" fill="#f2f2f2"/></g></svg>
        </g></g><g transform="translate(760 180)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_25" x1="9.01" y1="16.5" x2="9.01" y2="1.5" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#5e9641"/><stop offset=".34" stop-color="#6baa42"/><stop offset=".67" stop-color="#73b743"/><stop offset="1" stop-color="#76bb43"/></linearGradient></defs><title>Icon-networking-80</title><path d="M15.89 2.91h1.27a.34.34 0 0 1 .34.34v3.5a.34.34 0 0 1-.34.34h-1.27V2.91zm0 6.09h1.27a.34.34 0 0 1 .34.34v5.86a.34.34 0 0 1-.34.34h-1.27V9z" fill="#ffca00"/><rect x="2.13" y="1.5" width="13.76" height="15" rx=".69" fill="url(#ygc3_25)"/><path d="M5.9 12.9h-.71a.2.2 0 0 1-.19-.21V4.34a.19.19 0 0 1 .19-.2h1.93a.19.19 0 0 1 .19.2.2.2 0 0 1-.19.21H5.38v7.93h.52a.2.2 0 0 1 .19.21.21.21 0 0 1-.19.21z" fill="#b4ec36"/><path d="M6 13.92H4.4a.2.2 0 0 1-.19-.21L4.08 3.38a.2.2 0 0 1 .06-.15.16.16 0 0 1 .13-.06h2.85v.41H4.47l.12 9.92H6zm6-.92h-1.59a.19.19 0 0 1-.14-.07.18.18 0 0 1-.06-.14V7.9a.19.19 0 0 1 .19-.2h.91V5.45h.38v2.44a.2.2 0 0 1-.18.21h-.91v4.42H12z" fill="#b4ec36"/><rect x="7.07" y="2.29" width="6.14" height="3.11" rx=".26" fill="#365615"/><rect x="5.86" y="12.69" width="4.9" height="1.09" rx=".26" transform="rotate(90 8.305 13.235)" fill="#365615"/><rect x="3.99" y="12.71" width="4.9" height="1.09" rx=".26" transform="rotate(90 6.44 13.26)" fill="#365615"/><rect x="9.98" y="12.71" width="4.9" height="1.09" rx=".26" transform="rotate(90 12.425 13.255)" fill="#f2f2f2"/><ellipse cx="8.11" cy="8.06" rx="1.04" ry="1.12" fill="#f2f2f2"/><path d="M2.11 12.25H.84a.34.34 0 0 1-.34-.3V6.09a.34.34 0 0 1 .34-.34h1.27v6.5z" fill="#3b3b3b"/></g></svg>
        </g></g><g transform="translate(760 300)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_26" x1="8.88" y1="12.21" x2="8.88" y2=".21" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#0078d4"/><stop offset=".82" stop-color="#5ea0ef"/></linearGradient><linearGradient id="ygc3_27" x1="8.88" y1="16.84" x2="8.88" y2="12.21" gradientUnits="userSpaceOnUse"><stop offset=".15" stop-color="#ccc"/><stop offset="1" stop-color="#707070"/></linearGradient></defs><title>Icon-compute-21</title><rect x="-.12" y=".21" width="18" height="12" rx=".6" fill="url(#ygc3_26)"/><path fill="#50e6ff" d="M11.88 4.46v3.49l-3 1.76v-3.5l3-1.75z"/><path fill="#c3f1ff" d="M11.88 4.46l-3 1.76-3-1.76 3-1.75 3 1.75z"/><path fill="#9cebff" d="M8.88 6.22v3.49l-3-1.76V4.46l3 1.76z"/><path fill="#c3f1ff" d="M5.88 7.95l3-1.74v3.5l-3-1.76z"/><path fill="#9cebff" d="M11.88 7.95l-3-1.74v3.5l3-1.76z"/><path d="M12.49 15.84c-1.78-.28-1.85-1.56-1.85-3.63H7.11c0 2.07-.06 3.35-1.84 3.63a1 1 0 0 0-.89 1h9a1 1 0 0 0-.89-1z" fill="url(#ygc3_27)"/></g></svg>
        </g></g><g transform="translate(593.3333333333334 180)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_28" x1="9.01" y1="16.5" x2="9.01" y2="1.5" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#5e9641"/><stop offset=".34" stop-color="#6baa42"/><stop offset=".67" stop-color="#73b743"/><stop offset="1" stop-color="#76bb43"/></linearGradient></defs><title>Icon-networking-80</title><path d="M15.89 2.91h1.27a.34.34 0 0 1 .34.34v3.5a.34.34 0 0 1-.34.34h-1.27V2.91zm0 6.09h1.27a.34.34 0 0 1 .34.34v5.86a.34.34 0 0 1-.34.34h-1.27V9z" fill="#ffca00"/><rect x="2.13" y="1.5" width="13.76" height="15" rx=".69" fill="url(#ygc3_28)"/><path d="M5.9 12.9h-.71a.2.2 0 0 1-.19-.21V4.34a.19.19 0 0 1 .19-.2h1.93a.19.19 0 0 1 .19.2.2.2 0 0 1-.19.21H5.38v7.93h.52a.2.2 0 0 1 .19.21.21.21 0 0 1-.19.21z" fill="#b4ec36"/><path d="M6 13.92H4.4a.2.2 0 0 1-.19-.21L4.08 3.38a.2.2 0 0 1 .06-.15.16.16 0 0 1 .13-.06h2.85v.41H4.47l.12 9.92H6zm6-.92h-1.59a.19.19 0 0 1-.14-.07.18.18 0 0 1-.06-.14V7.9a.19.19 0 0 1 .19-.2h.91V5.45h.38v2.44a.2.2 0 0 1-.18.21h-.91v4.42H12z" fill="#b4ec36"/><rect x="7.07" y="2.29" width="6.14" height="3.11" rx=".26" fill="#365615"/><rect x="5.86" y="12.69" width="4.9" height="1.09" rx=".26" transform="rotate(90 8.305 13.235)" fill="#365615"/><rect x="3.99" y="12.71" width="4.9" height="1.09" rx=".26" transform="rotate(90 6.44 13.26)" fill="#365615"/><rect x="9.98" y="12.71" width="4.9" height="1.09" rx=".26" transform="rotate(90 12.425 13.255)" fill="#f2f2f2"/><ellipse cx="8.11" cy="8.06" rx="1.04" ry="1.12" fill="#f2f2f2"/><path d="M2.11 12.25H.84a.34.34 0 0 1-.34-.3V6.09a.34.34 0 0 1 .34-.34h1.27v6.5z" fill="#3b3b3b"/></g></svg>
        </g></g><g transform="translate(460 300)"><g transform="scale(2.78)">
            <svg svgBox="0 0 18 18" fill="msportalfx-svg-placeholder" role="presentation" focusable="false"><g><title/><defs><linearGradient id="ygc3_29" x1="8.88" y1="12.21" x2="8.88" y2=".21" gradientUnits="userSpaceOnUse"><stop offset="0" stop-color="#0078d4"/><stop offset=".82" stop-color="#5ea0ef"/></linearGradient><linearGradient id="ygc3_30" x1="8.88" y1="16.84" x2="8.88" y2="12.21" gradientUnits="userSpaceOnUse"><stop offset=".15" stop-color="#ccc"/><stop offset="1" stop-color="#707070"/></linearGradient></defs><title>Icon-compute-21</title><rect x="-.12" y=".21" width="18" height="12" rx=".6" fill="url(#ygc3_29)"/><path fill="#50e6ff" d="M11.88 4.46v3.49l-3 1.76v-3.5l3-1.75z"/><path fill="#c3f1ff" d="M11.88 4.46l-3 1.76-3-1.76 3-1.75 3 1.75z"/><path fill="#9cebff" d="M8.88 6.22v3.49l-3-1.76V4.46l3 1.76z"/><path fill="#c3f1ff" d="M5.88 7.95l3-1.74v3.5l-3-1.76z"/><path fill="#9cebff" d="M11.88 7.95l-3-1.74v3.5l3-1.76z"/><path d="M12.49 15.84c-1.78-.28-1.85-1.56-1.85-3.63H7.11c0 2.07-.06 3.35-1.84 3.63a1 1 0 0 0-.89 1h9a1 1 0 0 0-.89-1z" fill="url(#ygc3_30)"/></g></svg>
        </g></g><g transform="translate(155.64481051032817 46.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">ELK-VNET</text></g><g transform="translate(166.97652918901727 126.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">default</text></g><g transform="translate(148.63356605108754 226.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">elk-server394</text></g><g transform="translate(303.9740708189539 346.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">ELK-Server</text></g><g transform="translate(142.29647971292772 346.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">ELK-Server-nsg</text></g><g transform="translate(-2.697163457480727 346.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">ELK-Server-ip</text></g><g transform="translate(923.6594879545142 46.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">R_T</text></g><g transform="translate(916.9765291890172 126.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">default</text></g><g transform="translate(1329.9447304858206 226.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">jumpboxprovisione...</text></g><g transform="translate(1479.950592730352 346.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">JumpBoxProvisioner</text></g><g transform="translate(910.7596188637458 346.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">RT_NSG</text></g><g transform="translate(1326.9461924081438 346.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">JumpBoxProvisione...</text></g><g transform="translate(1061.9731034816912 226.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">web-326</text></g><g transform="translate(1210.7566877414802 346.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">Web-3-ip</text></g><g transform="translate(910.6335806063263 226.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">web1223</text></g><g transform="translate(1069.4269474030327 346.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">Web1</text></g><g transform="translate(597.2940431757225 346.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">RedTeamPool</text></g><g transform="translate(601.9662520670392 426.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">RedTeamLB</text></g><g transform="translate(605.7901301609555 516.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">RedTeamProbe</text></g><g transform="translate(441.43935554873053 516.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">LoadBalancerFront...</text></g><g transform="translate(760.6335806063263 226.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">web2790</text></g><g transform="translate(769.4269474030328 346.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">Web2</text></g><g transform="translate(593.9669139396597 226.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">web3796</text></g><g transform="translate(470.649225387775 346.578125)"><text font-family="Arial" font-size="12px" font-style="normal" font-weight="normal" text-anchor="start" fill="rgb(0,0,0)" fill-opacity="1" dy="1em" transform="translate(0 0)">web3</text></g></g></svg>
